module sevenseg (input [3:0] code, output [6:0]seg);

end module