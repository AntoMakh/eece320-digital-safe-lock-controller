module myModule();
    helapsojdjaoshda
endmodule