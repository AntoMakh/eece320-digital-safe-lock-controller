module myModule();
    
endmodule